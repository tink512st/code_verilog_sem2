`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/18/2025 08:10:24 PM
// Design Name: 
// Module Name: d_ff_posedge_posrst
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Reg_set(q1,q2,clk,rst,d1,d2);
input [7:0] d1,d2;
input clk,rst;
output reg [7:0] q1,q2;

always @(posedge clk ) begin
    if(rst) begin
        q1 <= 0;
        q2 <= 0;
     end
     else begin
        q1 <= d1;
        q2 <= d2;
     end
end
endmodule
