`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07/18/2025 09:50:20 PM
// Design Name: 
// Module Name: div_clk_to 40Hz
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module div_clk_t(clk,rst,clk_out,sel_an);
input [2:0] sel_an;
input clk,rst;
output reg clk_out;

parameter sys_freq = 100000000; //100Mhz
parameter count_scan = 50;

reg [7:0] slow_clk_freq; 
reg [21:0] K;
reg [20:0] counter;

always@(posedge clk) begin
    slow_clk_freq <= (count_scan * sel_an); 
    K <= sys_freq / slow_clk_freq;
end
always@(posedge clk, posedge rst) begin
    if(rst) begin
        counter <= 4'd1;
        clk_out <= 0;
    end
    else if(counter == K/2) begin
        clk_out <= ~clk_out;
        counter <= 1;
    end
    else 
        counter <= counter + 1;
end
endmodule
