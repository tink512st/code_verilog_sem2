module uartrx#(
	parameter clk_freq = 1000000, //1Mhz
	parameter baud_rate = 9600
)
(doneRx,rxData,clk,rst,rx);
input clk,rst;
input rx;
output reg doneRx;
output reg [7:0] rxData;

localparam clkcount = clk_freq/baud_rate;
reg [1:0] idle = 2'b00, start = 2'b01;
reg [1:0] state;

integer count = 0;
integer counts = 0;
reg uclk = 0;

always @(posedge clk) begin
	if(count < clkcount/2)
		count <= count + 1;
	else begin
		count <= 0;
		uclk <= ~uclk;
	end
end

always@(posedge uclk) begin
	if(rst) begin
		counts <= 0;
		doneRx <= 0;
		rxData <= 8'h00;
	end
	else begin
		case(state) 
			idle: begin
				counts <= 0;
				doneRx <= 0;
				rxData <= 8'h00;
				if(rx ==1'b0)
					state <= start;
				else 
					state <= idle;
			end
			start: begin
				if(counts<=7) begin
					rxData <= {rx,rxData[7:1]};
					counts <= counts + 1;
				end
				else begin
					counts <= 0;
					doneRx <= 1;
					state <= idle;
				end
			end
			default : state <= idle;
		endcase
	end
end
endmodule